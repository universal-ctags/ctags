module xyz

// static methods

enum Bosh {
    bim
    bam
}

fn Bosh.from_string(s string) !Bosh {
}

fn Bogus.nope() {
}
