module main
import os
import a.b.cd
