/*
*
**/
module top(outsig, insig);
output outsig;
input insig;
assign outsig = insig;
endmodule
