// #2738: processDesignElementL() go into infinite loop
interface static 0
