  // 6.16 String data type
  parameter string default_name = "John Smith"; // default_name:register => default_name:constant

  // 6.20 Constants
  parameter logic flag = 1 ; // flags:register => flags:constant
  parameter real r1 = 3.5e17; // r1:register => r1:constant
