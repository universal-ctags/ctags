// from UVM-1.2
`define defvar_with_comment \
  // comment in multi-line macro \
  logic foo;

`define defvar_without_comment \
  logic foo;
