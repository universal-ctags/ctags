function 0: