module aaa

enum Foo {
    aaa = 5
    bbb
    ccc
    @fn
    @struct
    ddd
}
