constant"	
