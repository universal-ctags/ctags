/* Legend:
 * <e> = empty (null)
 * <n> = non-empty
 */

module \ ;
	struct {
		struct {
			logic \ ;
			logic \eeen ;
		} \ ;
		struct {
			logic \ ;
			logic \eenn ;
		} \een ;
	} \ ;
	struct {
		struct {
			logic \ ;
			logic \enen ;
		} \ ;
		struct {
			logic \ ;
			logic \ennn ;
		} \enn ;
	} \en ;
endmodule

module \n ;
	struct {
		struct {
			logic \ ;
			logic \neen ;
		} \ ;
		struct {
			logic \ ;
			logic \nenn ;
		} \nen ;
	} \ ;
	struct {
		struct {
			logic \ ;
			logic \nnen ;
		} \ ;
		struct {
			logic \ ;
			logic \nnnn ;
		} \nnn ;
	} \nn ;
endmodule

