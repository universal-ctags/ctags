module xyz

fn (mut s Foo) yesnow() ! {
}
