module aaa

enum Foo {
    aaa = 5
    bbb
    ccc = C.foo
    @fn
    @struct [attr]
    ddd = 999  @[attr]
}
