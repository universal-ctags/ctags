-- https://www.ics.uci.edu/~jmoorkan/vhdlref/Synario%20VHDL%20Manual.pdf
entity logical_ops_1 is
  port (a, b, c, d: in bit;
        m: out bit);
end logical_ops_1;
