package body
