// Takne from #2413 submitted by @antoinemadec
typedef bit[31:0] int32_t;
module mod(
  input bit clk,
  input int32_t a
);
endmodule
